
module InstructionMem ( addrBus, dataBus );
  input [4:0] addrBus;
  output [7:0] dataBus;


endmodule

