
module DataMem_n8 ( AddrBus, Rd, Wr, LoadAcc, DataInBus, DataOutBus );
  input [4:0] AddrBus;
  input [7:0] DataInBus;
  output [7:0] DataOutBus;
  input Rd, Wr, LoadAcc;
  wire   N12, N13, N14, N15, N16, \DM[0][7] , \DM[0][6] , \DM[0][5] ,
         \DM[0][4] , \DM[0][3] , \DM[0][2] , \DM[0][1] , \DM[0][0] ,
         \DM[1][7] , \DM[1][6] , \DM[1][5] , \DM[1][4] , \DM[1][3] ,
         \DM[1][2] , \DM[1][1] , \DM[1][0] , \DM[2][7] , \DM[2][6] ,
         \DM[2][5] , \DM[2][4] , \DM[2][3] , \DM[2][2] , \DM[2][1] ,
         \DM[2][0] , \DM[3][7] , \DM[3][6] , \DM[3][5] , \DM[3][4] ,
         \DM[3][3] , \DM[3][2] , \DM[3][1] , \DM[3][0] , \DM[4][7] ,
         \DM[4][6] , \DM[4][5] , \DM[4][4] , \DM[4][3] , \DM[4][2] ,
         \DM[4][1] , \DM[4][0] , \DM[5][7] , \DM[5][6] , \DM[5][5] ,
         \DM[5][4] , \DM[5][3] , \DM[5][2] , \DM[5][1] , \DM[5][0] ,
         \DM[6][7] , \DM[6][6] , \DM[6][5] , \DM[6][4] , \DM[6][3] ,
         \DM[6][2] , \DM[6][1] , \DM[6][0] , \DM[7][7] , \DM[7][6] ,
         \DM[7][5] , \DM[7][4] , \DM[7][3] , \DM[7][2] , \DM[7][1] ,
         \DM[7][0] , \DM[8][7] , \DM[8][6] , \DM[8][5] , \DM[8][4] ,
         \DM[8][3] , \DM[8][2] , \DM[8][1] , \DM[8][0] , \DM[9][7] ,
         \DM[9][6] , \DM[9][5] , \DM[9][4] , \DM[9][3] , \DM[9][2] ,
         \DM[9][1] , \DM[9][0] , \DM[10][7] , \DM[10][6] , \DM[10][5] ,
         \DM[10][4] , \DM[10][3] , \DM[10][2] , \DM[10][1] , \DM[10][0] ,
         \DM[11][7] , \DM[11][6] , \DM[11][5] , \DM[11][4] , \DM[11][3] ,
         \DM[11][2] , \DM[11][1] , \DM[11][0] , \DM[12][7] , \DM[12][6] ,
         \DM[12][5] , \DM[12][4] , \DM[12][3] , \DM[12][2] , \DM[12][1] ,
         \DM[12][0] , \DM[13][7] , \DM[13][6] , \DM[13][5] , \DM[13][4] ,
         \DM[13][3] , \DM[13][2] , \DM[13][1] , \DM[13][0] , \DM[14][7] ,
         \DM[14][6] , \DM[14][5] , \DM[14][4] , \DM[14][3] , \DM[14][2] ,
         \DM[14][1] , \DM[14][0] , \DM[15][7] , \DM[15][6] , \DM[15][5] ,
         \DM[15][4] , \DM[15][3] , \DM[15][2] , \DM[15][1] , \DM[15][0] ,
         \DM[16][7] , \DM[16][6] , \DM[16][5] , \DM[16][4] , \DM[16][3] ,
         \DM[16][2] , \DM[16][1] , \DM[16][0] , \DM[17][7] , \DM[17][6] ,
         \DM[17][5] , \DM[17][4] , \DM[17][3] , \DM[17][2] , \DM[17][1] ,
         \DM[17][0] , \DM[18][7] , \DM[18][6] , \DM[18][5] , \DM[18][4] ,
         \DM[18][3] , \DM[18][2] , \DM[18][1] , \DM[18][0] , \DM[19][7] ,
         \DM[19][6] , \DM[19][5] , \DM[19][4] , \DM[19][3] , \DM[19][2] ,
         \DM[19][1] , \DM[19][0] , \DM[20][7] , \DM[20][6] , \DM[20][5] ,
         \DM[20][4] , \DM[20][3] , \DM[20][2] , \DM[20][1] , \DM[20][0] ,
         \DM[21][7] , \DM[21][6] , \DM[21][5] , \DM[21][4] , \DM[21][3] ,
         \DM[21][2] , \DM[21][1] , \DM[21][0] , \DM[22][7] , \DM[22][6] ,
         \DM[22][5] , \DM[22][4] , \DM[22][3] , \DM[22][2] , \DM[22][1] ,
         \DM[22][0] , \DM[23][7] , \DM[23][6] , \DM[23][5] , \DM[23][4] ,
         \DM[23][3] , \DM[23][2] , \DM[23][1] , \DM[23][0] , \DM[24][7] ,
         \DM[24][6] , \DM[24][5] , \DM[24][4] , \DM[24][3] , \DM[24][2] ,
         \DM[24][1] , \DM[24][0] , \DM[25][7] , \DM[25][6] , \DM[25][5] ,
         \DM[25][4] , \DM[25][3] , \DM[25][2] , \DM[25][1] , \DM[25][0] ,
         \DM[26][7] , \DM[26][6] , \DM[26][5] , \DM[26][4] , \DM[26][3] ,
         \DM[26][2] , \DM[26][1] , \DM[26][0] , \DM[27][7] , \DM[27][6] ,
         \DM[27][5] , \DM[27][4] , \DM[27][3] , \DM[27][2] , \DM[27][1] ,
         \DM[27][0] , \DM[28][7] , \DM[28][6] , \DM[28][5] , \DM[28][4] ,
         \DM[28][3] , \DM[28][2] , \DM[28][1] , \DM[28][0] , \DM[29][7] ,
         \DM[29][6] , \DM[29][5] , \DM[29][4] , \DM[29][3] , \DM[29][2] ,
         \DM[29][1] , \DM[29][0] , \DM[30][7] , \DM[30][6] , \DM[30][5] ,
         \DM[30][4] , \DM[30][3] , \DM[30][2] , \DM[30][1] , \DM[30][0] ,
         \DM[31][7] , \DM[31][6] , \DM[31][5] , \DM[31][4] , \DM[31][3] ,
         \DM[31][2] , \DM[31][1] , \DM[31][0] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153;
  assign N12 = AddrBus[0];
  assign N13 = AddrBus[1];
  assign N14 = AddrBus[2];
  assign N15 = AddrBus[3];
  assign N16 = AddrBus[4];

  LATCHX1 \DM_reg[0][7]  ( .CLK(n45), .D(DataInBus[7]), .Q(\DM[0][7] ) );
  LATCHX1 \DM_reg[0][6]  ( .CLK(n45), .D(DataInBus[6]), .Q(\DM[0][6] ) );
  LATCHX1 \DM_reg[0][5]  ( .CLK(n45), .D(DataInBus[5]), .Q(\DM[0][5] ) );
  LATCHX1 \DM_reg[0][4]  ( .CLK(n45), .D(DataInBus[4]), .Q(\DM[0][4] ) );
  LATCHX1 \DM_reg[0][3]  ( .CLK(n45), .D(DataInBus[3]), .Q(\DM[0][3] ) );
  LATCHX1 \DM_reg[0][2]  ( .CLK(n45), .D(DataInBus[2]), .Q(\DM[0][2] ) );
  LATCHX1 \DM_reg[0][1]  ( .CLK(n45), .D(DataInBus[1]), .Q(\DM[0][1] ) );
  LATCHX1 \DM_reg[0][0]  ( .CLK(n45), .D(DataInBus[0]), .Q(\DM[0][0] ) );
  LATCHX1 \DM_reg[1][7]  ( .CLK(n25), .D(DataInBus[7]), .Q(\DM[1][7] ) );
  LATCHX1 \DM_reg[1][6]  ( .CLK(n25), .D(DataInBus[6]), .Q(\DM[1][6] ) );
  LATCHX1 \DM_reg[1][5]  ( .CLK(n25), .D(DataInBus[5]), .Q(\DM[1][5] ) );
  LATCHX1 \DM_reg[1][4]  ( .CLK(n25), .D(DataInBus[4]), .Q(\DM[1][4] ) );
  LATCHX1 \DM_reg[1][3]  ( .CLK(n25), .D(DataInBus[3]), .Q(\DM[1][3] ) );
  LATCHX1 \DM_reg[1][2]  ( .CLK(n25), .D(DataInBus[2]), .Q(\DM[1][2] ) );
  LATCHX1 \DM_reg[1][1]  ( .CLK(n25), .D(DataInBus[1]), .Q(\DM[1][1] ) );
  LATCHX1 \DM_reg[1][0]  ( .CLK(n25), .D(DataInBus[0]), .Q(\DM[1][0] ) );
  LATCHX1 \DM_reg[2][7]  ( .CLK(n15), .D(DataInBus[7]), .Q(\DM[2][7] ) );
  LATCHX1 \DM_reg[2][6]  ( .CLK(n15), .D(DataInBus[6]), .Q(\DM[2][6] ) );
  LATCHX1 \DM_reg[2][5]  ( .CLK(n15), .D(DataInBus[5]), .Q(\DM[2][5] ) );
  LATCHX1 \DM_reg[2][4]  ( .CLK(n15), .D(DataInBus[4]), .Q(\DM[2][4] ) );
  LATCHX1 \DM_reg[2][3]  ( .CLK(n15), .D(DataInBus[3]), .Q(\DM[2][3] ) );
  LATCHX1 \DM_reg[2][2]  ( .CLK(n15), .D(DataInBus[2]), .Q(\DM[2][2] ) );
  LATCHX1 \DM_reg[2][1]  ( .CLK(n15), .D(DataInBus[1]), .Q(\DM[2][1] ) );
  LATCHX1 \DM_reg[2][0]  ( .CLK(n15), .D(DataInBus[0]), .Q(\DM[2][0] ) );
  LATCHX1 \DM_reg[3][7]  ( .CLK(n14), .D(DataInBus[7]), .Q(\DM[3][7] ) );
  LATCHX1 \DM_reg[3][6]  ( .CLK(n14), .D(DataInBus[6]), .Q(\DM[3][6] ) );
  LATCHX1 \DM_reg[3][5]  ( .CLK(n14), .D(DataInBus[5]), .Q(\DM[3][5] ) );
  LATCHX1 \DM_reg[3][4]  ( .CLK(n14), .D(DataInBus[4]), .Q(\DM[3][4] ) );
  LATCHX1 \DM_reg[3][3]  ( .CLK(n14), .D(DataInBus[3]), .Q(\DM[3][3] ) );
  LATCHX1 \DM_reg[3][2]  ( .CLK(n14), .D(DataInBus[2]), .Q(\DM[3][2] ) );
  LATCHX1 \DM_reg[3][1]  ( .CLK(n14), .D(DataInBus[1]), .Q(\DM[3][1] ) );
  LATCHX1 \DM_reg[3][0]  ( .CLK(n14), .D(DataInBus[0]), .Q(\DM[3][0] ) );
  LATCHX1 \DM_reg[4][7]  ( .CLK(n24), .D(DataInBus[7]), .Q(\DM[4][7] ) );
  LATCHX1 \DM_reg[4][6]  ( .CLK(n24), .D(DataInBus[6]), .Q(\DM[4][6] ) );
  LATCHX1 \DM_reg[4][5]  ( .CLK(n24), .D(DataInBus[5]), .Q(\DM[4][5] ) );
  LATCHX1 \DM_reg[4][4]  ( .CLK(n24), .D(DataInBus[4]), .Q(\DM[4][4] ) );
  LATCHX1 \DM_reg[4][3]  ( .CLK(n24), .D(DataInBus[3]), .Q(\DM[4][3] ) );
  LATCHX1 \DM_reg[4][2]  ( .CLK(n24), .D(DataInBus[2]), .Q(\DM[4][2] ) );
  LATCHX1 \DM_reg[4][1]  ( .CLK(n24), .D(DataInBus[1]), .Q(\DM[4][1] ) );
  LATCHX1 \DM_reg[4][0]  ( .CLK(n24), .D(DataInBus[0]), .Q(\DM[4][0] ) );
  LATCHX1 \DM_reg[5][7]  ( .CLK(n23), .D(DataInBus[7]), .Q(\DM[5][7] ) );
  LATCHX1 \DM_reg[5][6]  ( .CLK(n23), .D(DataInBus[6]), .Q(\DM[5][6] ) );
  LATCHX1 \DM_reg[5][5]  ( .CLK(n23), .D(DataInBus[5]), .Q(\DM[5][5] ) );
  LATCHX1 \DM_reg[5][4]  ( .CLK(n23), .D(DataInBus[4]), .Q(\DM[5][4] ) );
  LATCHX1 \DM_reg[5][3]  ( .CLK(n23), .D(DataInBus[3]), .Q(\DM[5][3] ) );
  LATCHX1 \DM_reg[5][2]  ( .CLK(n23), .D(DataInBus[2]), .Q(\DM[5][2] ) );
  LATCHX1 \DM_reg[5][1]  ( .CLK(n23), .D(DataInBus[1]), .Q(\DM[5][1] ) );
  LATCHX1 \DM_reg[5][0]  ( .CLK(n23), .D(DataInBus[0]), .Q(\DM[5][0] ) );
  LATCHX1 \DM_reg[6][7]  ( .CLK(n13), .D(DataInBus[7]), .Q(\DM[6][7] ) );
  LATCHX1 \DM_reg[6][6]  ( .CLK(n13), .D(DataInBus[6]), .Q(\DM[6][6] ) );
  LATCHX1 \DM_reg[6][5]  ( .CLK(n13), .D(DataInBus[5]), .Q(\DM[6][5] ) );
  LATCHX1 \DM_reg[6][4]  ( .CLK(n13), .D(DataInBus[4]), .Q(\DM[6][4] ) );
  LATCHX1 \DM_reg[6][3]  ( .CLK(n13), .D(DataInBus[3]), .Q(\DM[6][3] ) );
  LATCHX1 \DM_reg[6][2]  ( .CLK(n13), .D(DataInBus[2]), .Q(\DM[6][2] ) );
  LATCHX1 \DM_reg[6][1]  ( .CLK(n13), .D(DataInBus[1]), .Q(\DM[6][1] ) );
  LATCHX1 \DM_reg[6][0]  ( .CLK(n13), .D(DataInBus[0]), .Q(\DM[6][0] ) );
  LATCHX1 \DM_reg[7][7]  ( .CLK(n12), .D(DataInBus[7]), .Q(\DM[7][7] ) );
  LATCHX1 \DM_reg[7][6]  ( .CLK(n12), .D(DataInBus[6]), .Q(\DM[7][6] ) );
  LATCHX1 \DM_reg[7][5]  ( .CLK(n12), .D(DataInBus[5]), .Q(\DM[7][5] ) );
  LATCHX1 \DM_reg[7][4]  ( .CLK(n12), .D(DataInBus[4]), .Q(\DM[7][4] ) );
  LATCHX1 \DM_reg[7][3]  ( .CLK(n12), .D(DataInBus[3]), .Q(\DM[7][3] ) );
  LATCHX1 \DM_reg[7][2]  ( .CLK(n12), .D(DataInBus[2]), .Q(\DM[7][2] ) );
  LATCHX1 \DM_reg[7][1]  ( .CLK(n12), .D(DataInBus[1]), .Q(\DM[7][1] ) );
  LATCHX1 \DM_reg[7][0]  ( .CLK(n12), .D(DataInBus[0]), .Q(\DM[7][0] ) );
  LATCHX1 \DM_reg[8][7]  ( .CLK(n44), .D(DataInBus[7]), .Q(\DM[8][7] ) );
  LATCHX1 \DM_reg[8][6]  ( .CLK(n44), .D(DataInBus[6]), .Q(\DM[8][6] ) );
  LATCHX1 \DM_reg[8][5]  ( .CLK(n44), .D(DataInBus[5]), .Q(\DM[8][5] ) );
  LATCHX1 \DM_reg[8][4]  ( .CLK(n44), .D(DataInBus[4]), .Q(\DM[8][4] ) );
  LATCHX1 \DM_reg[8][3]  ( .CLK(n44), .D(DataInBus[3]), .Q(\DM[8][3] ) );
  LATCHX1 \DM_reg[8][2]  ( .CLK(n44), .D(DataInBus[2]), .Q(\DM[8][2] ) );
  LATCHX1 \DM_reg[8][1]  ( .CLK(n44), .D(DataInBus[1]), .Q(\DM[8][1] ) );
  LATCHX1 \DM_reg[8][0]  ( .CLK(n44), .D(DataInBus[0]), .Q(\DM[8][0] ) );
  LATCHX1 \DM_reg[9][7]  ( .CLK(n22), .D(DataInBus[7]), .Q(\DM[9][7] ) );
  LATCHX1 \DM_reg[9][6]  ( .CLK(n22), .D(DataInBus[6]), .Q(\DM[9][6] ) );
  LATCHX1 \DM_reg[9][5]  ( .CLK(n22), .D(DataInBus[5]), .Q(\DM[9][5] ) );
  LATCHX1 \DM_reg[9][4]  ( .CLK(n22), .D(DataInBus[4]), .Q(\DM[9][4] ) );
  LATCHX1 \DM_reg[9][3]  ( .CLK(n22), .D(DataInBus[3]), .Q(\DM[9][3] ) );
  LATCHX1 \DM_reg[9][2]  ( .CLK(n22), .D(DataInBus[2]), .Q(\DM[9][2] ) );
  LATCHX1 \DM_reg[9][1]  ( .CLK(n22), .D(DataInBus[1]), .Q(\DM[9][1] ) );
  LATCHX1 \DM_reg[9][0]  ( .CLK(n22), .D(DataInBus[0]), .Q(\DM[9][0] ) );
  LATCHX1 \DM_reg[10][7]  ( .CLK(n11), .D(DataInBus[7]), .Q(\DM[10][7] ) );
  LATCHX1 \DM_reg[10][6]  ( .CLK(n11), .D(DataInBus[6]), .Q(\DM[10][6] ) );
  LATCHX1 \DM_reg[10][5]  ( .CLK(n11), .D(DataInBus[5]), .Q(\DM[10][5] ) );
  LATCHX1 \DM_reg[10][4]  ( .CLK(n11), .D(DataInBus[4]), .Q(\DM[10][4] ) );
  LATCHX1 \DM_reg[10][3]  ( .CLK(n11), .D(DataInBus[3]), .Q(\DM[10][3] ) );
  LATCHX1 \DM_reg[10][2]  ( .CLK(n11), .D(DataInBus[2]), .Q(\DM[10][2] ) );
  LATCHX1 \DM_reg[10][1]  ( .CLK(n11), .D(DataInBus[1]), .Q(\DM[10][1] ) );
  LATCHX1 \DM_reg[10][0]  ( .CLK(n11), .D(DataInBus[0]), .Q(\DM[10][0] ) );
  LATCHX1 \DM_reg[11][7]  ( .CLK(n10), .D(DataInBus[7]), .Q(\DM[11][7] ) );
  LATCHX1 \DM_reg[11][6]  ( .CLK(n10), .D(DataInBus[6]), .Q(\DM[11][6] ) );
  LATCHX1 \DM_reg[11][5]  ( .CLK(n10), .D(DataInBus[5]), .Q(\DM[11][5] ) );
  LATCHX1 \DM_reg[11][4]  ( .CLK(n10), .D(DataInBus[4]), .Q(\DM[11][4] ) );
  LATCHX1 \DM_reg[11][3]  ( .CLK(n10), .D(DataInBus[3]), .Q(\DM[11][3] ) );
  LATCHX1 \DM_reg[11][2]  ( .CLK(n10), .D(DataInBus[2]), .Q(\DM[11][2] ) );
  LATCHX1 \DM_reg[11][1]  ( .CLK(n10), .D(DataInBus[1]), .Q(\DM[11][1] ) );
  LATCHX1 \DM_reg[11][0]  ( .CLK(n10), .D(DataInBus[0]), .Q(\DM[11][0] ) );
  LATCHX1 \DM_reg[12][7]  ( .CLK(n21), .D(DataInBus[7]), .Q(\DM[12][7] ) );
  LATCHX1 \DM_reg[12][6]  ( .CLK(n21), .D(DataInBus[6]), .Q(\DM[12][6] ) );
  LATCHX1 \DM_reg[12][5]  ( .CLK(n21), .D(DataInBus[5]), .Q(\DM[12][5] ) );
  LATCHX1 \DM_reg[12][4]  ( .CLK(n21), .D(DataInBus[4]), .Q(\DM[12][4] ) );
  LATCHX1 \DM_reg[12][3]  ( .CLK(n21), .D(DataInBus[3]), .Q(\DM[12][3] ) );
  LATCHX1 \DM_reg[12][2]  ( .CLK(n21), .D(DataInBus[2]), .Q(\DM[12][2] ) );
  LATCHX1 \DM_reg[12][1]  ( .CLK(n21), .D(DataInBus[1]), .Q(\DM[12][1] ) );
  LATCHX1 \DM_reg[12][0]  ( .CLK(n21), .D(DataInBus[0]), .Q(\DM[12][0] ) );
  LATCHX1 \DM_reg[13][7]  ( .CLK(n20), .D(DataInBus[7]), .Q(\DM[13][7] ) );
  LATCHX1 \DM_reg[13][6]  ( .CLK(n20), .D(DataInBus[6]), .Q(\DM[13][6] ) );
  LATCHX1 \DM_reg[13][5]  ( .CLK(n20), .D(DataInBus[5]), .Q(\DM[13][5] ) );
  LATCHX1 \DM_reg[13][4]  ( .CLK(n20), .D(DataInBus[4]), .Q(\DM[13][4] ) );
  LATCHX1 \DM_reg[13][3]  ( .CLK(n20), .D(DataInBus[3]), .Q(\DM[13][3] ) );
  LATCHX1 \DM_reg[13][2]  ( .CLK(n20), .D(DataInBus[2]), .Q(\DM[13][2] ) );
  LATCHX1 \DM_reg[13][1]  ( .CLK(n20), .D(DataInBus[1]), .Q(\DM[13][1] ) );
  LATCHX1 \DM_reg[13][0]  ( .CLK(n20), .D(DataInBus[0]), .Q(\DM[13][0] ) );
  LATCHX1 \DM_reg[14][7]  ( .CLK(n9), .D(DataInBus[7]), .Q(\DM[14][7] ) );
  LATCHX1 \DM_reg[14][6]  ( .CLK(n9), .D(DataInBus[6]), .Q(\DM[14][6] ) );
  LATCHX1 \DM_reg[14][5]  ( .CLK(n9), .D(DataInBus[5]), .Q(\DM[14][5] ) );
  LATCHX1 \DM_reg[14][4]  ( .CLK(n9), .D(DataInBus[4]), .Q(\DM[14][4] ) );
  LATCHX1 \DM_reg[14][3]  ( .CLK(n9), .D(DataInBus[3]), .Q(\DM[14][3] ) );
  LATCHX1 \DM_reg[14][2]  ( .CLK(n9), .D(DataInBus[2]), .Q(\DM[14][2] ) );
  LATCHX1 \DM_reg[14][1]  ( .CLK(n9), .D(DataInBus[1]), .Q(\DM[14][1] ) );
  LATCHX1 \DM_reg[14][0]  ( .CLK(n9), .D(DataInBus[0]), .Q(\DM[14][0] ) );
  LATCHX1 \DM_reg[15][7]  ( .CLK(n8), .D(DataInBus[7]), .Q(\DM[15][7] ) );
  LATCHX1 \DM_reg[15][6]  ( .CLK(n8), .D(DataInBus[6]), .Q(\DM[15][6] ) );
  LATCHX1 \DM_reg[15][5]  ( .CLK(n8), .D(DataInBus[5]), .Q(\DM[15][5] ) );
  LATCHX1 \DM_reg[15][4]  ( .CLK(n8), .D(DataInBus[4]), .Q(\DM[15][4] ) );
  LATCHX1 \DM_reg[15][3]  ( .CLK(n8), .D(DataInBus[3]), .Q(\DM[15][3] ) );
  LATCHX1 \DM_reg[15][2]  ( .CLK(n8), .D(DataInBus[2]), .Q(\DM[15][2] ) );
  LATCHX1 \DM_reg[15][1]  ( .CLK(n8), .D(DataInBus[1]), .Q(\DM[15][1] ) );
  LATCHX1 \DM_reg[15][0]  ( .CLK(n8), .D(DataInBus[0]), .Q(\DM[15][0] ) );
  LATCHX1 \DM_reg[16][7]  ( .CLK(n35), .D(DataInBus[7]), .Q(\DM[16][7] ) );
  LATCHX1 \DM_reg[16][6]  ( .CLK(n35), .D(DataInBus[6]), .Q(\DM[16][6] ) );
  LATCHX1 \DM_reg[16][5]  ( .CLK(n35), .D(DataInBus[5]), .Q(\DM[16][5] ) );
  LATCHX1 \DM_reg[16][4]  ( .CLK(n35), .D(DataInBus[4]), .Q(\DM[16][4] ) );
  LATCHX1 \DM_reg[16][3]  ( .CLK(n35), .D(DataInBus[3]), .Q(\DM[16][3] ) );
  LATCHX1 \DM_reg[16][2]  ( .CLK(n35), .D(DataInBus[2]), .Q(\DM[16][2] ) );
  LATCHX1 \DM_reg[16][1]  ( .CLK(n35), .D(DataInBus[1]), .Q(\DM[16][1] ) );
  LATCHX1 \DM_reg[16][0]  ( .CLK(n35), .D(DataInBus[0]), .Q(\DM[16][0] ) );
  LATCHX1 \DM_reg[17][7]  ( .CLK(n34), .D(DataInBus[7]), .Q(\DM[17][7] ) );
  LATCHX1 \DM_reg[17][6]  ( .CLK(n34), .D(DataInBus[6]), .Q(\DM[17][6] ) );
  LATCHX1 \DM_reg[17][5]  ( .CLK(n34), .D(DataInBus[5]), .Q(\DM[17][5] ) );
  LATCHX1 \DM_reg[17][4]  ( .CLK(n34), .D(DataInBus[4]), .Q(\DM[17][4] ) );
  LATCHX1 \DM_reg[17][3]  ( .CLK(n34), .D(DataInBus[3]), .Q(\DM[17][3] ) );
  LATCHX1 \DM_reg[17][2]  ( .CLK(n34), .D(DataInBus[2]), .Q(\DM[17][2] ) );
  LATCHX1 \DM_reg[17][1]  ( .CLK(n34), .D(DataInBus[1]), .Q(\DM[17][1] ) );
  LATCHX1 \DM_reg[17][0]  ( .CLK(n34), .D(DataInBus[0]), .Q(\DM[17][0] ) );
  LATCHX1 \DM_reg[18][7]  ( .CLK(n33), .D(DataInBus[7]), .Q(\DM[18][7] ) );
  LATCHX1 \DM_reg[18][6]  ( .CLK(n33), .D(DataInBus[6]), .Q(\DM[18][6] ) );
  LATCHX1 \DM_reg[18][5]  ( .CLK(n33), .D(DataInBus[5]), .Q(\DM[18][5] ) );
  LATCHX1 \DM_reg[18][4]  ( .CLK(n33), .D(DataInBus[4]), .Q(\DM[18][4] ) );
  LATCHX1 \DM_reg[18][3]  ( .CLK(n33), .D(DataInBus[3]), .Q(\DM[18][3] ) );
  LATCHX1 \DM_reg[18][2]  ( .CLK(n33), .D(DataInBus[2]), .Q(\DM[18][2] ) );
  LATCHX1 \DM_reg[18][1]  ( .CLK(n33), .D(DataInBus[1]), .Q(\DM[18][1] ) );
  LATCHX1 \DM_reg[18][0]  ( .CLK(n33), .D(DataInBus[0]), .Q(\DM[18][0] ) );
  LATCHX1 \DM_reg[19][7]  ( .CLK(n32), .D(DataInBus[7]), .Q(\DM[19][7] ) );
  LATCHX1 \DM_reg[19][6]  ( .CLK(n32), .D(DataInBus[6]), .Q(\DM[19][6] ) );
  LATCHX1 \DM_reg[19][5]  ( .CLK(n32), .D(DataInBus[5]), .Q(\DM[19][5] ) );
  LATCHX1 \DM_reg[19][4]  ( .CLK(n32), .D(DataInBus[4]), .Q(\DM[19][4] ) );
  LATCHX1 \DM_reg[19][3]  ( .CLK(n32), .D(DataInBus[3]), .Q(\DM[19][3] ) );
  LATCHX1 \DM_reg[19][2]  ( .CLK(n32), .D(DataInBus[2]), .Q(\DM[19][2] ) );
  LATCHX1 \DM_reg[19][1]  ( .CLK(n32), .D(DataInBus[1]), .Q(\DM[19][1] ) );
  LATCHX1 \DM_reg[19][0]  ( .CLK(n32), .D(DataInBus[0]), .Q(\DM[19][0] ) );
  LATCHX1 \DM_reg[20][7]  ( .CLK(n31), .D(DataInBus[7]), .Q(\DM[20][7] ) );
  LATCHX1 \DM_reg[20][6]  ( .CLK(n31), .D(DataInBus[6]), .Q(\DM[20][6] ) );
  LATCHX1 \DM_reg[20][5]  ( .CLK(n31), .D(DataInBus[5]), .Q(\DM[20][5] ) );
  LATCHX1 \DM_reg[20][4]  ( .CLK(n31), .D(DataInBus[4]), .Q(\DM[20][4] ) );
  LATCHX1 \DM_reg[20][3]  ( .CLK(n31), .D(DataInBus[3]), .Q(\DM[20][3] ) );
  LATCHX1 \DM_reg[20][2]  ( .CLK(n31), .D(DataInBus[2]), .Q(\DM[20][2] ) );
  LATCHX1 \DM_reg[20][1]  ( .CLK(n31), .D(DataInBus[1]), .Q(\DM[20][1] ) );
  LATCHX1 \DM_reg[20][0]  ( .CLK(n31), .D(DataInBus[0]), .Q(\DM[20][0] ) );
  LATCHX1 \DM_reg[21][7]  ( .CLK(n30), .D(DataInBus[7]), .Q(\DM[21][7] ) );
  LATCHX1 \DM_reg[21][6]  ( .CLK(n30), .D(DataInBus[6]), .Q(\DM[21][6] ) );
  LATCHX1 \DM_reg[21][5]  ( .CLK(n30), .D(DataInBus[5]), .Q(\DM[21][5] ) );
  LATCHX1 \DM_reg[21][4]  ( .CLK(n30), .D(DataInBus[4]), .Q(\DM[21][4] ) );
  LATCHX1 \DM_reg[21][3]  ( .CLK(n30), .D(DataInBus[3]), .Q(\DM[21][3] ) );
  LATCHX1 \DM_reg[21][2]  ( .CLK(n30), .D(DataInBus[2]), .Q(\DM[21][2] ) );
  LATCHX1 \DM_reg[21][1]  ( .CLK(n30), .D(DataInBus[1]), .Q(\DM[21][1] ) );
  LATCHX1 \DM_reg[21][0]  ( .CLK(n30), .D(DataInBus[0]), .Q(\DM[21][0] ) );
  LATCHX1 \DM_reg[22][7]  ( .CLK(n29), .D(DataInBus[7]), .Q(\DM[22][7] ) );
  LATCHX1 \DM_reg[22][6]  ( .CLK(n29), .D(DataInBus[6]), .Q(\DM[22][6] ) );
  LATCHX1 \DM_reg[22][5]  ( .CLK(n29), .D(DataInBus[5]), .Q(\DM[22][5] ) );
  LATCHX1 \DM_reg[22][4]  ( .CLK(n29), .D(DataInBus[4]), .Q(\DM[22][4] ) );
  LATCHX1 \DM_reg[22][3]  ( .CLK(n29), .D(DataInBus[3]), .Q(\DM[22][3] ) );
  LATCHX1 \DM_reg[22][2]  ( .CLK(n29), .D(DataInBus[2]), .Q(\DM[22][2] ) );
  LATCHX1 \DM_reg[22][1]  ( .CLK(n29), .D(DataInBus[1]), .Q(\DM[22][1] ) );
  LATCHX1 \DM_reg[22][0]  ( .CLK(n29), .D(DataInBus[0]), .Q(\DM[22][0] ) );
  LATCHX1 \DM_reg[23][7]  ( .CLK(n28), .D(DataInBus[7]), .Q(\DM[23][7] ) );
  LATCHX1 \DM_reg[23][6]  ( .CLK(n28), .D(DataInBus[6]), .Q(\DM[23][6] ) );
  LATCHX1 \DM_reg[23][5]  ( .CLK(n28), .D(DataInBus[5]), .Q(\DM[23][5] ) );
  LATCHX1 \DM_reg[23][4]  ( .CLK(n28), .D(DataInBus[4]), .Q(\DM[23][4] ) );
  LATCHX1 \DM_reg[23][3]  ( .CLK(n28), .D(DataInBus[3]), .Q(\DM[23][3] ) );
  LATCHX1 \DM_reg[23][2]  ( .CLK(n28), .D(DataInBus[2]), .Q(\DM[23][2] ) );
  LATCHX1 \DM_reg[23][1]  ( .CLK(n28), .D(DataInBus[1]), .Q(\DM[23][1] ) );
  LATCHX1 \DM_reg[23][0]  ( .CLK(n28), .D(DataInBus[0]), .Q(\DM[23][0] ) );
  LATCHX1 \DM_reg[24][7]  ( .CLK(n43), .D(DataInBus[7]), .Q(\DM[24][7] ) );
  LATCHX1 \DM_reg[24][6]  ( .CLK(n43), .D(DataInBus[6]), .Q(\DM[24][6] ) );
  LATCHX1 \DM_reg[24][5]  ( .CLK(n43), .D(DataInBus[5]), .Q(\DM[24][5] ) );
  LATCHX1 \DM_reg[24][4]  ( .CLK(n43), .D(DataInBus[4]), .Q(\DM[24][4] ) );
  LATCHX1 \DM_reg[24][3]  ( .CLK(n43), .D(DataInBus[3]), .Q(\DM[24][3] ) );
  LATCHX1 \DM_reg[24][2]  ( .CLK(n43), .D(DataInBus[2]), .Q(\DM[24][2] ) );
  LATCHX1 \DM_reg[24][1]  ( .CLK(n43), .D(DataInBus[1]), .Q(\DM[24][1] ) );
  LATCHX1 \DM_reg[24][0]  ( .CLK(n43), .D(DataInBus[0]), .Q(\DM[24][0] ) );
  LATCHX1 \DM_reg[25][7]  ( .CLK(n42), .D(DataInBus[7]), .Q(\DM[25][7] ) );
  LATCHX1 \DM_reg[25][6]  ( .CLK(n42), .D(DataInBus[6]), .Q(\DM[25][6] ) );
  LATCHX1 \DM_reg[25][5]  ( .CLK(n42), .D(DataInBus[5]), .Q(\DM[25][5] ) );
  LATCHX1 \DM_reg[25][4]  ( .CLK(n42), .D(DataInBus[4]), .Q(\DM[25][4] ) );
  LATCHX1 \DM_reg[25][3]  ( .CLK(n42), .D(DataInBus[3]), .Q(\DM[25][3] ) );
  LATCHX1 \DM_reg[25][2]  ( .CLK(n42), .D(DataInBus[2]), .Q(\DM[25][2] ) );
  LATCHX1 \DM_reg[25][1]  ( .CLK(n42), .D(DataInBus[1]), .Q(\DM[25][1] ) );
  LATCHX1 \DM_reg[25][0]  ( .CLK(n42), .D(DataInBus[0]), .Q(\DM[25][0] ) );
  LATCHX1 \DM_reg[26][7]  ( .CLK(n41), .D(DataInBus[7]), .Q(\DM[26][7] ) );
  LATCHX1 \DM_reg[26][6]  ( .CLK(n41), .D(DataInBus[6]), .Q(\DM[26][6] ) );
  LATCHX1 \DM_reg[26][5]  ( .CLK(n41), .D(DataInBus[5]), .Q(\DM[26][5] ) );
  LATCHX1 \DM_reg[26][4]  ( .CLK(n41), .D(DataInBus[4]), .Q(\DM[26][4] ) );
  LATCHX1 \DM_reg[26][3]  ( .CLK(n41), .D(DataInBus[3]), .Q(\DM[26][3] ) );
  LATCHX1 \DM_reg[26][2]  ( .CLK(n41), .D(DataInBus[2]), .Q(\DM[26][2] ) );
  LATCHX1 \DM_reg[26][1]  ( .CLK(n41), .D(DataInBus[1]), .Q(\DM[26][1] ) );
  LATCHX1 \DM_reg[26][0]  ( .CLK(n41), .D(DataInBus[0]), .Q(\DM[26][0] ) );
  LATCHX1 \DM_reg[27][7]  ( .CLK(n40), .D(DataInBus[7]), .Q(\DM[27][7] ) );
  LATCHX1 \DM_reg[27][6]  ( .CLK(n40), .D(DataInBus[6]), .Q(\DM[27][6] ) );
  LATCHX1 \DM_reg[27][5]  ( .CLK(n40), .D(DataInBus[5]), .Q(\DM[27][5] ) );
  LATCHX1 \DM_reg[27][4]  ( .CLK(n40), .D(DataInBus[4]), .Q(\DM[27][4] ) );
  LATCHX1 \DM_reg[27][3]  ( .CLK(n40), .D(DataInBus[3]), .Q(\DM[27][3] ) );
  LATCHX1 \DM_reg[27][2]  ( .CLK(n40), .D(DataInBus[2]), .Q(\DM[27][2] ) );
  LATCHX1 \DM_reg[27][1]  ( .CLK(n40), .D(DataInBus[1]), .Q(\DM[27][1] ) );
  LATCHX1 \DM_reg[27][0]  ( .CLK(n40), .D(DataInBus[0]), .Q(\DM[27][0] ) );
  LATCHX1 \DM_reg[28][7]  ( .CLK(n39), .D(DataInBus[7]), .Q(\DM[28][7] ) );
  LATCHX1 \DM_reg[28][6]  ( .CLK(n39), .D(DataInBus[6]), .Q(\DM[28][6] ) );
  LATCHX1 \DM_reg[28][5]  ( .CLK(n39), .D(DataInBus[5]), .Q(\DM[28][5] ) );
  LATCHX1 \DM_reg[28][4]  ( .CLK(n39), .D(DataInBus[4]), .Q(\DM[28][4] ) );
  LATCHX1 \DM_reg[28][3]  ( .CLK(n39), .D(DataInBus[3]), .Q(\DM[28][3] ) );
  LATCHX1 \DM_reg[28][2]  ( .CLK(n39), .D(DataInBus[2]), .Q(\DM[28][2] ) );
  LATCHX1 \DM_reg[28][1]  ( .CLK(n39), .D(DataInBus[1]), .Q(\DM[28][1] ) );
  LATCHX1 \DM_reg[28][0]  ( .CLK(n39), .D(DataInBus[0]), .Q(\DM[28][0] ) );
  LATCHX1 \DM_reg[29][7]  ( .CLK(n38), .D(DataInBus[7]), .Q(\DM[29][7] ) );
  LATCHX1 \DM_reg[29][6]  ( .CLK(n38), .D(DataInBus[6]), .Q(\DM[29][6] ) );
  LATCHX1 \DM_reg[29][5]  ( .CLK(n38), .D(DataInBus[5]), .Q(\DM[29][5] ) );
  LATCHX1 \DM_reg[29][4]  ( .CLK(n38), .D(DataInBus[4]), .Q(\DM[29][4] ) );
  LATCHX1 \DM_reg[29][3]  ( .CLK(n38), .D(DataInBus[3]), .Q(\DM[29][3] ) );
  LATCHX1 \DM_reg[29][2]  ( .CLK(n38), .D(DataInBus[2]), .Q(\DM[29][2] ) );
  LATCHX1 \DM_reg[29][1]  ( .CLK(n38), .D(DataInBus[1]), .Q(\DM[29][1] ) );
  LATCHX1 \DM_reg[29][0]  ( .CLK(n38), .D(DataInBus[0]), .Q(\DM[29][0] ) );
  LATCHX1 \DM_reg[30][7]  ( .CLK(n37), .D(DataInBus[7]), .Q(\DM[30][7] ) );
  LATCHX1 \DM_reg[30][6]  ( .CLK(n37), .D(DataInBus[6]), .Q(\DM[30][6] ) );
  LATCHX1 \DM_reg[30][5]  ( .CLK(n37), .D(DataInBus[5]), .Q(\DM[30][5] ) );
  LATCHX1 \DM_reg[30][4]  ( .CLK(n37), .D(DataInBus[4]), .Q(\DM[30][4] ) );
  LATCHX1 \DM_reg[30][3]  ( .CLK(n37), .D(DataInBus[3]), .Q(\DM[30][3] ) );
  LATCHX1 \DM_reg[30][2]  ( .CLK(n37), .D(DataInBus[2]), .Q(\DM[30][2] ) );
  LATCHX1 \DM_reg[30][1]  ( .CLK(n37), .D(DataInBus[1]), .Q(\DM[30][1] ) );
  LATCHX1 \DM_reg[30][0]  ( .CLK(n37), .D(DataInBus[0]), .Q(\DM[30][0] ) );
  LATCHX1 \DM_reg[31][7]  ( .CLK(n36), .D(DataInBus[7]), .Q(\DM[31][7] ) );
  LATCHX1 \DM_reg[31][6]  ( .CLK(n36), .D(DataInBus[6]), .Q(\DM[31][6] ) );
  LATCHX1 \DM_reg[31][5]  ( .CLK(n36), .D(DataInBus[5]), .Q(\DM[31][5] ) );
  LATCHX1 \DM_reg[31][4]  ( .CLK(n36), .D(DataInBus[4]), .Q(\DM[31][4] ) );
  LATCHX1 \DM_reg[31][3]  ( .CLK(n36), .D(DataInBus[3]), .Q(\DM[31][3] ) );
  LATCHX1 \DM_reg[31][2]  ( .CLK(n36), .D(DataInBus[2]), .Q(\DM[31][2] ) );
  LATCHX1 \DM_reg[31][1]  ( .CLK(n36), .D(DataInBus[1]), .Q(\DM[31][1] ) );
  LATCHX1 \DM_reg[31][0]  ( .CLK(n36), .D(DataInBus[0]), .Q(\DM[31][0] ) );
  MUX41X1 U2 ( .IN1(\DM[4][7] ), .IN3(\DM[6][7] ), .IN2(\DM[5][7] ), .IN4(
        \DM[7][7] ), .S0(n5), .S1(n58), .Q(n141) );
  MUX41X1 U3 ( .IN1(\DM[0][7] ), .IN3(\DM[2][7] ), .IN2(\DM[1][7] ), .IN4(
        \DM[3][7] ), .S0(n5), .S1(n56), .Q(n143) );
  MUX41X1 U4 ( .IN1(\DM[8][7] ), .IN3(\DM[10][7] ), .IN2(\DM[9][7] ), .IN4(
        \DM[11][7] ), .S0(n61), .S1(n57), .Q(n142) );
  MUX41X1 U5 ( .IN1(\DM[12][7] ), .IN3(\DM[14][7] ), .IN2(\DM[13][7] ), .IN4(
        \DM[15][7] ), .S0(n61), .S1(n1), .Q(n140) );
  MUX41X1 U6 ( .IN1(\DM[16][7] ), .IN3(\DM[18][7] ), .IN2(\DM[17][7] ), .IN4(
        \DM[19][7] ), .S0(n5), .S1(n59), .Q(n147) );
  MUX41X1 U7 ( .IN1(\DM[24][7] ), .IN3(\DM[26][7] ), .IN2(\DM[25][7] ), .IN4(
        \DM[27][7] ), .S0(n5), .S1(n2), .Q(n146) );
  MUX41X1 U8 ( .IN1(\DM[28][7] ), .IN3(\DM[30][7] ), .IN2(\DM[29][7] ), .IN4(
        \DM[31][7] ), .S0(n5), .S1(n2), .Q(n144) );
  MUX41X1 U9 ( .IN1(\DM[20][7] ), .IN3(\DM[22][7] ), .IN2(\DM[21][7] ), .IN4(
        \DM[23][7] ), .S0(n5), .S1(n1), .Q(n145) );
  MUX41X1 U10 ( .IN1(\DM[28][6] ), .IN3(\DM[30][6] ), .IN2(\DM[29][6] ), .IN4(
        \DM[31][6] ), .S0(n61), .S1(n58), .Q(n133) );
  MUX41X1 U11 ( .IN1(\DM[24][6] ), .IN3(\DM[26][6] ), .IN2(\DM[25][6] ), .IN4(
        \DM[27][6] ), .S0(n5), .S1(n56), .Q(n135) );
  MUX41X1 U12 ( .IN1(\DM[20][6] ), .IN3(\DM[22][6] ), .IN2(\DM[21][6] ), .IN4(
        \DM[23][6] ), .S0(n5), .S1(n57), .Q(n134) );
  AND3X1 U13 ( .IN1(n7), .IN2(n151), .IN3(n59), .Q(n50) );
  AND3X1 U14 ( .IN1(n7), .IN2(n151), .IN3(n60), .Q(n51) );
  IBUFFX4 U15 ( .INP(n60), .ZN(n57) );
  INVX0 U16 ( .INP(N13), .ZN(n3) );
  IBUFFX4 U17 ( .INP(n60), .ZN(n56) );
  MUX41X1 U18 ( .IN1(n66), .IN3(n64), .IN2(n65), .IN4(n63), .S0(N14), .S1(N12), 
        .Q(n72) );
  MUX41X1 U19 ( .IN1(\DM[7][0] ), .IN3(\DM[5][0] ), .IN2(\DM[15][0] ), .IN4(
        \DM[13][0] ), .S0(n6), .S1(N15), .Q(n63) );
  MUX41X1 U20 ( .IN1(\DM[26][0] ), .IN3(\DM[24][0] ), .IN2(\DM[27][0] ), .IN4(
        \DM[25][0] ), .S0(n6), .S1(N12), .Q(n69) );
  IBUFFX4 U21 ( .INP(n60), .ZN(n1) );
  IBUFFX16 U22 ( .INP(n60), .ZN(n2) );
  IBUFFX16 U23 ( .INP(n60), .ZN(n59) );
  MUX21X1 U24 ( .IN1(n72), .IN2(n71), .S(N16), .Q(n73) );
  MUX41X1 U25 ( .IN1(\DM[6][0] ), .IN3(\DM[4][0] ), .IN2(\DM[14][0] ), .IN4(
        \DM[12][0] ), .S0(n6), .S1(N15), .Q(n64) );
  NBUFFX2 U26 ( .INP(N13), .Z(n4) );
  IBUFFX4 U27 ( .INP(n3), .ZN(n61) );
  IBUFFX4 U28 ( .INP(n3), .ZN(n5) );
  INVX0 U29 ( .INP(N13), .ZN(n6) );
  INVX0 U30 ( .INP(n61), .ZN(n7) );
  IBUFFX4 U31 ( .INP(N12), .ZN(n60) );
  AND2X1 U32 ( .IN1(n16), .IN2(n26), .Q(n8) );
  AND2X1 U33 ( .IN1(n16), .IN2(n19), .Q(n9) );
  AND2X1 U34 ( .IN1(n16), .IN2(n27), .Q(n10) );
  AND2X1 U35 ( .IN1(n16), .IN2(n18), .Q(n11) );
  AND2X1 U36 ( .IN1(n17), .IN2(n26), .Q(n12) );
  AND2X1 U37 ( .IN1(n17), .IN2(n19), .Q(n13) );
  AND2X1 U38 ( .IN1(n17), .IN2(n27), .Q(n14) );
  AND2X1 U39 ( .IN1(n17), .IN2(n18), .Q(n15) );
  INVX0 U40 ( .INP(n55), .ZN(n152) );
  INVX2 U41 ( .INP(n60), .ZN(n58) );
  AND3X1 U42 ( .IN1(Wr), .IN2(n153), .IN3(n55), .Q(n16) );
  AND3X1 U43 ( .IN1(n152), .IN2(n153), .IN3(Wr), .Q(n17) );
  AND3X1 U44 ( .IN1(n60), .IN2(n151), .IN3(n61), .Q(n18) );
  AND3X1 U45 ( .IN1(n61), .IN2(n60), .IN3(n52), .Q(n19) );
  AND2X1 U46 ( .IN1(n16), .IN2(n48), .Q(n20) );
  AND2X1 U47 ( .IN1(n16), .IN2(n49), .Q(n21) );
  AND2X1 U48 ( .IN1(n16), .IN2(n50), .Q(n22) );
  AND2X1 U49 ( .IN1(n17), .IN2(n48), .Q(n23) );
  AND2X1 U50 ( .IN1(n17), .IN2(n49), .Q(n24) );
  AND2X1 U51 ( .IN1(n17), .IN2(n50), .Q(n25) );
  AND3X1 U52 ( .IN1(n61), .IN2(n59), .IN3(n54), .Q(n26) );
  AND3X1 U53 ( .IN1(n59), .IN2(n151), .IN3(n61), .Q(n27) );
  AND2X1 U54 ( .IN1(n26), .IN2(n46), .Q(n28) );
  AND2X1 U55 ( .IN1(n19), .IN2(n46), .Q(n29) );
  AND2X1 U56 ( .IN1(n48), .IN2(n46), .Q(n30) );
  AND2X1 U57 ( .IN1(n49), .IN2(n46), .Q(n31) );
  AND2X1 U58 ( .IN1(n27), .IN2(n46), .Q(n32) );
  AND2X1 U59 ( .IN1(n18), .IN2(n46), .Q(n33) );
  AND2X1 U60 ( .IN1(n50), .IN2(n46), .Q(n34) );
  AND2X1 U61 ( .IN1(n51), .IN2(n46), .Q(n35) );
  AND2X1 U62 ( .IN1(n26), .IN2(n47), .Q(n36) );
  AND2X1 U63 ( .IN1(n19), .IN2(n47), .Q(n37) );
  AND2X1 U64 ( .IN1(n48), .IN2(n47), .Q(n38) );
  AND2X1 U65 ( .IN1(n49), .IN2(n47), .Q(n39) );
  AND2X1 U66 ( .IN1(n27), .IN2(n47), .Q(n40) );
  AND2X1 U67 ( .IN1(n18), .IN2(n47), .Q(n41) );
  AND2X1 U68 ( .IN1(n50), .IN2(n47), .Q(n42) );
  AND2X1 U69 ( .IN1(n51), .IN2(n47), .Q(n43) );
  AND2X1 U70 ( .IN1(n51), .IN2(n16), .Q(n44) );
  AND2X1 U71 ( .IN1(n51), .IN2(n17), .Q(n45) );
  INVX0 U72 ( .INP(n53), .ZN(n151) );
  INVX0 U73 ( .INP(n3), .ZN(n62) );
  NBUFFX2 U74 ( .INP(N14), .Z(n52) );
  NBUFFX2 U75 ( .INP(N14), .Z(n53) );
  NBUFFX2 U76 ( .INP(N14), .Z(n54) );
  AND3X1 U77 ( .IN1(Wr), .IN2(n152), .IN3(N16), .Q(n46) );
  AND3X1 U78 ( .IN1(n55), .IN2(Wr), .IN3(N16), .Q(n47) );
  AND3X1 U79 ( .IN1(n59), .IN2(n7), .IN3(n53), .Q(n48) );
  AND3X1 U80 ( .IN1(n60), .IN2(n7), .IN3(n54), .Q(n49) );
  MUX21X1 U81 ( .IN1(\DM[0][3] ), .IN2(n106), .S(Rd), .Q(DataOutBus[3]) );
  MUX21X1 U82 ( .IN1(\DM[0][4] ), .IN2(n117), .S(Rd), .Q(DataOutBus[4]) );
  MUX21X1 U83 ( .IN1(\DM[0][6] ), .IN2(n139), .S(Rd), .Q(DataOutBus[6]) );
  MUX21X1 U84 ( .IN1(\DM[0][7] ), .IN2(n150), .S(Rd), .Q(DataOutBus[7]) );
  NBUFFX2 U85 ( .INP(N15), .Z(n55) );
  INVX0 U86 ( .INP(N16), .ZN(n153) );
  MUX41X1 U87 ( .IN1(\DM[0][0] ), .IN3(\DM[2][0] ), .IN2(\DM[8][0] ), .IN4(
        \DM[10][0] ), .S0(n4), .S1(N15), .Q(n66) );
  MUX41X1 U88 ( .IN1(\DM[1][0] ), .IN3(\DM[3][0] ), .IN2(\DM[9][0] ), .IN4(
        \DM[11][0] ), .S0(n62), .S1(N15), .Q(n65) );
  MUX41X1 U89 ( .IN1(\DM[16][0] ), .IN3(\DM[18][0] ), .IN2(\DM[17][0] ), .IN4(
        \DM[19][0] ), .S0(n4), .S1(N12), .Q(n70) );
  MUX41X1 U90 ( .IN1(\DM[20][0] ), .IN3(\DM[22][0] ), .IN2(\DM[21][0] ), .IN4(
        \DM[23][0] ), .S0(n4), .S1(N12), .Q(n68) );
  MUX41X1 U91 ( .IN1(\DM[28][0] ), .IN3(\DM[30][0] ), .IN2(\DM[29][0] ), .IN4(
        \DM[31][0] ), .S0(n4), .S1(N12), .Q(n67) );
  MUX41X1 U92 ( .IN1(n70), .IN3(n69), .IN2(n68), .IN4(n67), .S0(n55), .S1(n53), 
        .Q(n71) );
  MUX21X1 U93 ( .IN1(\DM[0][0] ), .IN2(n73), .S(Rd), .Q(DataOutBus[0]) );
  MUX41X1 U94 ( .IN1(\DM[0][1] ), .IN3(\DM[2][1] ), .IN2(\DM[1][1] ), .IN4(
        \DM[3][1] ), .S0(n61), .S1(n58), .Q(n77) );
  MUX41X1 U95 ( .IN1(\DM[8][1] ), .IN3(\DM[10][1] ), .IN2(\DM[9][1] ), .IN4(
        \DM[11][1] ), .S0(n61), .S1(n59), .Q(n76) );
  MUX41X1 U96 ( .IN1(\DM[4][1] ), .IN3(\DM[6][1] ), .IN2(\DM[5][1] ), .IN4(
        \DM[7][1] ), .S0(n61), .S1(n2), .Q(n75) );
  MUX41X1 U97 ( .IN1(\DM[12][1] ), .IN3(\DM[14][1] ), .IN2(\DM[13][1] ), .IN4(
        \DM[15][1] ), .S0(n5), .S1(n56), .Q(n74) );
  MUX41X1 U98 ( .IN1(n77), .IN3(n76), .IN2(n75), .IN4(n74), .S0(n55), .S1(n54), 
        .Q(n83) );
  MUX41X1 U99 ( .IN1(\DM[16][1] ), .IN3(\DM[18][1] ), .IN2(\DM[17][1] ), .IN4(
        \DM[19][1] ), .S0(n4), .S1(n1), .Q(n81) );
  MUX41X1 U100 ( .IN1(\DM[24][1] ), .IN3(\DM[26][1] ), .IN2(\DM[25][1] ), 
        .IN4(\DM[27][1] ), .S0(n4), .S1(n56), .Q(n80) );
  MUX41X1 U101 ( .IN1(\DM[20][1] ), .IN3(\DM[22][1] ), .IN2(\DM[21][1] ), 
        .IN4(\DM[23][1] ), .S0(n4), .S1(n57), .Q(n79) );
  MUX41X1 U102 ( .IN1(\DM[28][1] ), .IN3(\DM[30][1] ), .IN2(\DM[29][1] ), 
        .IN4(\DM[31][1] ), .S0(n5), .S1(n1), .Q(n78) );
  MUX41X1 U103 ( .IN1(n81), .IN3(n80), .IN2(n79), .IN4(n78), .S0(n55), .S1(n52), .Q(n82) );
  MUX21X1 U104 ( .IN1(n83), .IN2(n82), .S(N16), .Q(n84) );
  MUX21X1 U105 ( .IN1(\DM[0][1] ), .IN2(n84), .S(Rd), .Q(DataOutBus[1]) );
  MUX41X1 U106 ( .IN1(\DM[0][2] ), .IN3(\DM[2][2] ), .IN2(\DM[1][2] ), .IN4(
        \DM[3][2] ), .S0(n61), .S1(n2), .Q(n88) );
  MUX41X1 U107 ( .IN1(\DM[8][2] ), .IN3(\DM[10][2] ), .IN2(\DM[9][2] ), .IN4(
        \DM[11][2] ), .S0(n61), .S1(n1), .Q(n87) );
  MUX41X1 U108 ( .IN1(\DM[4][2] ), .IN3(\DM[6][2] ), .IN2(\DM[5][2] ), .IN4(
        \DM[7][2] ), .S0(n5), .S1(n56), .Q(n86) );
  MUX41X1 U109 ( .IN1(\DM[12][2] ), .IN3(\DM[14][2] ), .IN2(\DM[13][2] ), 
        .IN4(\DM[15][2] ), .S0(n61), .S1(n58), .Q(n85) );
  MUX41X1 U110 ( .IN1(n88), .IN3(n87), .IN2(n86), .IN4(n85), .S0(n55), .S1(n53), .Q(n94) );
  MUX41X1 U111 ( .IN1(\DM[16][2] ), .IN3(\DM[18][2] ), .IN2(\DM[17][2] ), 
        .IN4(\DM[19][2] ), .S0(n5), .S1(n57), .Q(n92) );
  MUX41X1 U112 ( .IN1(\DM[24][2] ), .IN3(\DM[26][2] ), .IN2(\DM[25][2] ), 
        .IN4(\DM[27][2] ), .S0(n61), .S1(n58), .Q(n91) );
  MUX41X1 U113 ( .IN1(\DM[20][2] ), .IN3(\DM[22][2] ), .IN2(\DM[21][2] ), 
        .IN4(\DM[23][2] ), .S0(n61), .S1(n59), .Q(n90) );
  MUX41X1 U114 ( .IN1(\DM[28][2] ), .IN3(\DM[30][2] ), .IN2(\DM[29][2] ), 
        .IN4(\DM[31][2] ), .S0(n5), .S1(n57), .Q(n89) );
  MUX41X1 U115 ( .IN1(n92), .IN3(n91), .IN2(n90), .IN4(n89), .S0(n55), .S1(n54), .Q(n93) );
  MUX21X1 U116 ( .IN1(n94), .IN2(n93), .S(N16), .Q(n95) );
  MUX21X1 U117 ( .IN1(\DM[0][2] ), .IN2(n95), .S(Rd), .Q(DataOutBus[2]) );
  MUX41X1 U118 ( .IN1(\DM[0][3] ), .IN3(\DM[2][3] ), .IN2(\DM[1][3] ), .IN4(
        \DM[3][3] ), .S0(n61), .S1(n56), .Q(n99) );
  MUX41X1 U119 ( .IN1(\DM[8][3] ), .IN3(\DM[10][3] ), .IN2(\DM[9][3] ), .IN4(
        \DM[11][3] ), .S0(n5), .S1(n57), .Q(n98) );
  MUX41X1 U120 ( .IN1(\DM[4][3] ), .IN3(\DM[6][3] ), .IN2(\DM[5][3] ), .IN4(
        \DM[7][3] ), .S0(n61), .S1(n58), .Q(n97) );
  MUX41X1 U121 ( .IN1(\DM[12][3] ), .IN3(\DM[14][3] ), .IN2(\DM[13][3] ), 
        .IN4(\DM[15][3] ), .S0(n61), .S1(n2), .Q(n96) );
  MUX41X1 U122 ( .IN1(n99), .IN3(n98), .IN2(n97), .IN4(n96), .S0(n55), .S1(n52), .Q(n105) );
  MUX41X1 U123 ( .IN1(\DM[16][3] ), .IN3(\DM[18][3] ), .IN2(\DM[17][3] ), 
        .IN4(\DM[19][3] ), .S0(n5), .S1(n59), .Q(n103) );
  MUX41X1 U124 ( .IN1(\DM[24][3] ), .IN3(\DM[26][3] ), .IN2(\DM[25][3] ), 
        .IN4(\DM[27][3] ), .S0(n61), .S1(n2), .Q(n102) );
  MUX41X1 U125 ( .IN1(\DM[20][3] ), .IN3(\DM[22][3] ), .IN2(\DM[21][3] ), 
        .IN4(\DM[23][3] ), .S0(n5), .S1(n1), .Q(n101) );
  MUX41X1 U126 ( .IN1(\DM[28][3] ), .IN3(\DM[30][3] ), .IN2(\DM[29][3] ), 
        .IN4(\DM[31][3] ), .S0(n5), .S1(n59), .Q(n100) );
  MUX41X1 U127 ( .IN1(n103), .IN3(n102), .IN2(n101), .IN4(n100), .S0(n55), 
        .S1(n53), .Q(n104) );
  MUX21X1 U128 ( .IN1(n105), .IN2(n104), .S(N16), .Q(n106) );
  MUX41X1 U129 ( .IN1(\DM[0][4] ), .IN3(\DM[2][4] ), .IN2(\DM[1][4] ), .IN4(
        \DM[3][4] ), .S0(n61), .S1(n58), .Q(n110) );
  MUX41X1 U130 ( .IN1(\DM[8][4] ), .IN3(\DM[10][4] ), .IN2(\DM[9][4] ), .IN4(
        \DM[11][4] ), .S0(n5), .S1(n59), .Q(n109) );
  MUX41X1 U131 ( .IN1(\DM[4][4] ), .IN3(\DM[6][4] ), .IN2(\DM[5][4] ), .IN4(
        \DM[7][4] ), .S0(n61), .S1(n2), .Q(n108) );
  MUX41X1 U132 ( .IN1(\DM[12][4] ), .IN3(\DM[14][4] ), .IN2(\DM[13][4] ), 
        .IN4(\DM[15][4] ), .S0(n61), .S1(n56), .Q(n107) );
  MUX41X1 U133 ( .IN1(n110), .IN3(n109), .IN2(n108), .IN4(n107), .S0(n55), 
        .S1(n54), .Q(n116) );
  MUX41X1 U134 ( .IN1(\DM[16][4] ), .IN3(\DM[18][4] ), .IN2(\DM[17][4] ), 
        .IN4(\DM[19][4] ), .S0(n61), .S1(n1), .Q(n114) );
  MUX41X1 U135 ( .IN1(\DM[24][4] ), .IN3(\DM[26][4] ), .IN2(\DM[25][4] ), 
        .IN4(\DM[27][4] ), .S0(n5), .S1(n56), .Q(n113) );
  MUX41X1 U136 ( .IN1(\DM[20][4] ), .IN3(\DM[22][4] ), .IN2(\DM[21][4] ), 
        .IN4(\DM[23][4] ), .S0(n61), .S1(n57), .Q(n112) );
  MUX41X1 U137 ( .IN1(\DM[28][4] ), .IN3(\DM[30][4] ), .IN2(\DM[29][4] ), 
        .IN4(\DM[31][4] ), .S0(n5), .S1(n1), .Q(n111) );
  MUX41X1 U138 ( .IN1(n114), .IN3(n113), .IN2(n112), .IN4(n111), .S0(n55), 
        .S1(n52), .Q(n115) );
  MUX21X1 U139 ( .IN1(n116), .IN2(n115), .S(N16), .Q(n117) );
  MUX41X1 U140 ( .IN1(\DM[0][5] ), .IN3(\DM[2][5] ), .IN2(\DM[1][5] ), .IN4(
        \DM[3][5] ), .S0(n61), .S1(n2), .Q(n121) );
  MUX41X1 U141 ( .IN1(\DM[8][5] ), .IN3(\DM[10][5] ), .IN2(\DM[9][5] ), .IN4(
        \DM[11][5] ), .S0(n61), .S1(n1), .Q(n120) );
  MUX41X1 U142 ( .IN1(\DM[4][5] ), .IN3(\DM[6][5] ), .IN2(\DM[5][5] ), .IN4(
        \DM[7][5] ), .S0(n5), .S1(n56), .Q(n119) );
  MUX41X1 U143 ( .IN1(\DM[12][5] ), .IN3(\DM[14][5] ), .IN2(\DM[13][5] ), 
        .IN4(\DM[15][5] ), .S0(n5), .S1(n58), .Q(n118) );
  MUX41X1 U144 ( .IN1(n121), .IN3(n120), .IN2(n119), .IN4(n118), .S0(n55), 
        .S1(n53), .Q(n127) );
  MUX41X1 U145 ( .IN1(\DM[16][5] ), .IN3(\DM[18][5] ), .IN2(\DM[17][5] ), 
        .IN4(\DM[19][5] ), .S0(n61), .S1(n57), .Q(n125) );
  MUX41X1 U146 ( .IN1(\DM[24][5] ), .IN3(\DM[26][5] ), .IN2(\DM[25][5] ), 
        .IN4(\DM[27][5] ), .S0(n5), .S1(n58), .Q(n124) );
  MUX41X1 U147 ( .IN1(\DM[20][5] ), .IN3(\DM[22][5] ), .IN2(\DM[21][5] ), 
        .IN4(\DM[23][5] ), .S0(n5), .S1(n59), .Q(n123) );
  MUX41X1 U148 ( .IN1(\DM[28][5] ), .IN3(\DM[30][5] ), .IN2(\DM[29][5] ), 
        .IN4(\DM[31][5] ), .S0(n61), .S1(n57), .Q(n122) );
  MUX41X1 U149 ( .IN1(n125), .IN3(n124), .IN2(n123), .IN4(n122), .S0(n55), 
        .S1(n54), .Q(n126) );
  MUX21X1 U150 ( .IN1(n127), .IN2(n126), .S(N16), .Q(n128) );
  MUX21X1 U151 ( .IN1(\DM[0][5] ), .IN2(n128), .S(Rd), .Q(DataOutBus[5]) );
  MUX41X1 U152 ( .IN1(\DM[0][6] ), .IN3(\DM[2][6] ), .IN2(\DM[1][6] ), .IN4(
        \DM[3][6] ), .S0(n5), .S1(n1), .Q(n132) );
  MUX41X1 U153 ( .IN1(\DM[8][6] ), .IN3(\DM[10][6] ), .IN2(\DM[9][6] ), .IN4(
        \DM[11][6] ), .S0(n5), .S1(n56), .Q(n131) );
  MUX41X1 U154 ( .IN1(\DM[4][6] ), .IN3(\DM[6][6] ), .IN2(\DM[5][6] ), .IN4(
        \DM[7][6] ), .S0(n61), .S1(n57), .Q(n130) );
  MUX41X1 U155 ( .IN1(\DM[12][6] ), .IN3(\DM[14][6] ), .IN2(\DM[13][6] ), 
        .IN4(\DM[15][6] ), .S0(n5), .S1(n58), .Q(n129) );
  MUX41X1 U156 ( .IN1(n132), .IN3(n131), .IN2(n130), .IN4(n129), .S0(n55), 
        .S1(n52), .Q(n138) );
  MUX41X1 U157 ( .IN1(\DM[16][6] ), .IN3(\DM[18][6] ), .IN2(\DM[17][6] ), 
        .IN4(\DM[19][6] ), .S0(n5), .S1(n2), .Q(n136) );
  MUX41X1 U158 ( .IN1(n136), .IN3(n135), .IN2(n134), .IN4(n133), .S0(n55), 
        .S1(n53), .Q(n137) );
  MUX21X1 U159 ( .IN1(n138), .IN2(n137), .S(N16), .Q(n139) );
  MUX41X1 U160 ( .IN1(n143), .IN3(n142), .IN2(n141), .IN4(n140), .S0(n55), 
        .S1(n54), .Q(n149) );
  MUX41X1 U161 ( .IN1(n147), .IN3(n146), .IN2(n145), .IN4(n144), .S0(n55), 
        .S1(n52), .Q(n148) );
  MUX21X1 U162 ( .IN1(n149), .IN2(n148), .S(N16), .Q(n150) );
endmodule

